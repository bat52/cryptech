
`ifdef DUMP_EN
dump localdump();
`endif